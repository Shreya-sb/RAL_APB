`include "interface.sv"
`include "reg_block.sv"
`include "seq_item.sv"
`include "adapter.sv"
`include "reg_seq.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
