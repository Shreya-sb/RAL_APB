`include "reg_block.sv"
`include "reg_seq.sv"
`include "adapter.sv"
`include "registers.sv"
`include "seq_item.sv"
`include "sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "environment.sv"
`include "interface.sv"
